//module multiplexer_4_1
//(
//	input input0,
//	input input1,
//	input input2,
//	input input3,
//	input [1:0] sel,
//	output reg out
//);
//	always @(*)
//	begin
//		
//	end